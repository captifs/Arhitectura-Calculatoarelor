module hello_world(
    output out,
    input in
    );
 
    not(out, in);
 
endmodule
